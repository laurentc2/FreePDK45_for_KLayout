* INV circuit for Double inverter LVS check

.SUBCKT INV A Z gnd vdd
M1 gnd A Z gnd NMOS_GVT L=0.05U W=0.095U
M2 vdd A Z vdd PMOS_GVT L=0.05U W=0.27U
.ENDS INV

.SUBCKT DBLE_INV_SPLIT A ZA ZB gnd vdd
X1 A ZA gnd vdd INV
X1 A ZB gnd vdd INV
.ENDS DBLE_INV_SPLIT

.SUBCKT DBLE_INV_MERGE A ZA ZB gnd vdd
X1 A ZA gnd vdd INV
X1 A ZB gnd vdd INV
.ENDS DBLE_INV_MERGE